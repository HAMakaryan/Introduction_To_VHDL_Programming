LIBRARY IEEE;                   -- IEEE library
USE IEEE.STD_LOGIC_1164.ALL;    -- Necessary to use the std_logic

ENTITY my_circuit_name IS
  PORT(
    inp1  : IN  STD_LOGIC;    --Input  port
    inp2  : IN  STD_LOGIC;    --Input  port
    outp1 : OUT STD_LOGIC;    --Output port
    outp2 : OUT STD_LOGIC;    --Output port
    outp3 : OUT STD_LOGIC     --Output port
  );
END my_circuit_name;





